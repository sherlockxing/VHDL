NET "I_sys_clk_50M" TNM_NET = I_sys_clk_50M;
TIMESPEC TS_I_sys_clk_50M = PERIOD "I_sys_clk_50M" 20 ns HIGH 50%;

NET "I_sys_clk_50M"    LOC = Y6       |   IOSTANDARD = LVCMOS33;  
NET I_sys_rst_50M        LOC = U5       |   IOSTANDARD = LVCMOS33; 
NET I_start                      LOC = R6     |   IOSTANDARD = LVCMOS33;
NET I_stop                      LOC = T6    |   IOSTANDARD = LVCMOS33;   
#NET O_row0_en             LOC = V7       |  IOSTANDARD = LVCMOS33;  
NET "led_dout[0]"     LOC = U22     |  IOSTANDARD = LVCMOS33;  
NET "led_dout[1]"     LOC = T22      |  IOSTANDARD = LVCMOS33;
NET "led_dout[2]"     LOC = W20    |  IOSTANDARD = LVCMOS33;
NET "led_dout[3]"     LOC = W21    |  IOSTANDARD = LVCMOS33;
NET "led_dout[4]"     LOC = U20     |  IOSTANDARD = LVCMOS33; 
NET "led_dout[5]"     LOC = U21     |  IOSTANDARD = LVCMOS33;  
NET "led_dout[6]"     LOC = W22    |  IOSTANDARD = LVCMOS33;
NET "led_dout[7]"     LOC = V22     |  IOSTANDARD = LVCMOS33;
NET "I_sys_rst_50M" CLOCK_DEDICATED_ROUTE = FALSE;

